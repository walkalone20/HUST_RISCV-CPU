`define PROG_PATH(name) `"C:/Users/Desktop/cpu21-riscv/programs/name.hex`"
